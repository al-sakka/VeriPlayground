-- Hello There this is a normal comment
-- Hello There this is a normal comment
